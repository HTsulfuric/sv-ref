package wide_pkg;
    typedef struct packed {
        logic [63:0] upper;
        logic [63:0] lower;
    } wide128_t;
endpackage
