package test_pkg;
    typedef struct packed {
        logic signed [7:0] signed_val;
        logic [7:0] unsigned_val;
    } mixed_t;
endpackage
